library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity generato_sin_wave is 
port ( clk:in std_logic ;
dataout : out integer  range  -128 to 127);
end generato_sin_wave;
architecture behavioral of generato_sin_wave is 
signal i : integer range 0 to 29:=0;
type type_memory is array (0 to 29) of integer range -128 to 127;
type memory_type is array (0 to 29) of integer range -128 to 127;
--ROM for storing the sine values generated by MATLAB.
signal sine : memory_type :=(0,16,31,45,58,67,74,77,77,74,67,58,45,31,16,0,
-16,-31,-45,-58,-67,-74,-77,-77,-74,-67,-58,-45,-31,-16);

begin

process(clk)
begin
  --to check the rising edge of the clock signal
if(rising_edge(clk)) then    
dataout <= sine(i);
i <= i+ 1;
if(i = 29) then
i <= 0;
end if;
end if;
end process;

end Behavioral;


